<?xml version="1.0" encoding="utf-8" standalone="no" ?> <svg version="1.0" xmlns="http://www.w3.org/2000/svg"> <g fill="#000000" stroke="none"> <path d="M3600 12374 c-221 -15 -362 -27 -465 -40 -729 -91 -1321 -315 -1780 -675 -119 -93 -317 -292 -396 -399 -170 -229 -275 -472 -331 -770 -19 -96 -22 -152 -23 -340 0 -194 3 -240 22 -335 40 -195 103 -355 196 -499 217 -332 548 -535 960 -586 125 -16 403 -7 507 15 251 55 448 162 633 343 199 195 311 432 339 714 44 454 -160 879 -612 1273 -123 107 -150 141 -142 180 13 72 170 179 342 235 213 69 530 77 790 20 124 -26 201 -54 325 -115 401 -198 708 -627 855 -1194 134 -515 154 -1238 49 -1766 -84 -423 -249 -765 -483 -1001 -158 -160 -310 -248 -515 -301 -130 -33 -263 -39 -514 -22 -117 8 -289 14 -382 14 l-170 0 -67 -33 c-77 -38 -171 -127 -211 -200 -124 -228 -36 -500 198 -612 127 -61 284 -73 590 -45 206 19 303 19 433 -1 268 -40 476 -145 668 -338 261 -264 438 -668 529 -1210 36 -217 53 -395 67 -693 24 -529 -26 -1002 -143 -1369 -218 -681 -644 -1103 -1237 -1223 -222 -46 -505 -52 -712 -16 -309 54 -618 230 -662 378 l-12 39 50 47 c28 25 105 92 172 149 299 253 484 542 553 862 29 137 32 389 6 523 -80 404 -343 718 -737 880 -192 79 -378 111 -645 111 -215 0 -305 -12 -472 -60 -345 -99 -672 -375 -839 -707 -135 -268 -181 -623 -127 -982 85 -573 421 -1063 1005 -1468 614 -426 1386 -656 2293 -686 1451 -47 2614 329 3380 1094 423 422 662 897 756 1505 20 125 23 185 23 440 1 312 -6 399 -50 650 -220 1232 -1121 2032 -2739 2431 -110 27 -208 49 -217 49 -42 0 -12 17 70 39 48 13 190 57 316 98 1174 382 1881 924 2201 1688 125 298 174 554 182 943 7 369 -15 584 -93 881 -47 182 -91 297 -184 486 -162 328 -384 604 -676 839 -526 423 -1180 662 -2029 742 -150 14 -724 26 -845 18z"/> </g> </svg>