<svg version="1.0">

<g
fill="#000000" stroke="none">
<path d="M4495 12298 c-604 -535 -1486 -866 -2660 -998 -331 -37 -854 -70
-1104 -70 l-101 0 -2 -415 -3 -416 30 -29 30 -29 735 -4 c620 -3 753 -7 850
-21 149 -22 254 -50 316 -86 82 -46 123 -142 161 -372 16 -95 18 -371 21
-3663 2 -2593 0 -3591 -8 -3675 -44 -446 -177 -714 -416 -838 -279 -144 -663
-202 -1350 -202 l-330 0 -27 -28 -27 -28 0 -389 0 -389 27 -28 27 -28 3386 0
3386 0 27 28 27 28 0 390 0 390 -27 26 -28 26 -390 5 c-415 5 -557 17 -779 62
-212 43 -367 103 -480 187 -156 115 -260 347 -312 693 -17 114 -18 350 -21
5005 l-3 4884 -27 28 -27 28 -410 -1 -411 0 -80 -71z"/>
</g>
</svg>
